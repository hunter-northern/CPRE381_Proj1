
library IEEE;
use IEEE.std_logic_1164.all;

entity decoder5t32 is

  port(i_S  : in std_logic_vector (4 downto 0);
	o_Y : out std_logic_vector(31 downto 0));

end decoder5t32;

architecture structure of decoder5t32 is
begin

o_Y <=
"00000000000000000000000000000001" when i_S = "00000" else
"00000000000000000000000000000010" when i_S = "00001" else
"00000000000000000000000000000100" when i_S = "00010" else
"00000000000000000000000000001000" when i_S = "00011" else
"00000000000000000000000000010000" when i_S = "00100" else
"00000000000000000000000000100000" when i_S = "00101" else
"00000000000000000000000001000000" when i_S = "00110" else
"00000000000000000000000010000000" when i_S = "00111" else
"00000000000000000000000100000000" when i_S = "01000" else
"00000000000000000000001000000000" when i_S = "01001" else
"00000000000000000000010000000000" when i_S = "01010" else
"00000000000000000000100000000000" when i_S = "01011" else
"00000000000000000001000000000000" when i_S = "01100" else
"00000000000000000010000000000000" when i_S = "01101" else
"00000000000000000100000000000000" when i_S = "01110" else
"00000000000000001000000000000000" when i_S = "01111" else
"00000000000000010000000000000000" when i_S = "10000" else
"00000000000000100000000000000000" when i_S = "10001" else
"00000000000001000000000000000000" when i_S = "10010" else
"00000000000010000000000000000000" when i_S = "10011" else
"00000000000100000000000000000000" when i_S = "10100" else
"00000000001000000000000000000000" when i_S = "10101" else
"00000000010000000000000000000000" when i_S = "10110" else
"00000000100000000000000000000000" when i_S = "10111" else
"00000001000000000000000000000000" when i_S = "11000" else
"00000010000000000000000000000000" when i_S = "11001" else
"00000100000000000000000000000000" when i_S = "11010" else
"00001000000000000000000000000000" when i_S = "11011" else
"00010000000000000000000000000000" when i_S = "11100" else
"00100000000000000000000000000000" when i_S = "11101" else
"01000000000000000000000000000000" when i_S = "11110" else
"10000000000000000000000000000000" when i_S = "11111" else
"00000000000000000000000000000000";
end structure;